`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   19:40:34 06/28/2016
// Design Name:   main
// Module Name:   F:/ali/home work/verilog/project/project2/test4.v
// Project Name:  project2
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: main
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module test4;

	// Inputs
	reg clk;

	// Instantiate the Unit Under Test (UUT)
	main uut (
		.clk(clk)
	);

	initial begin
		// Initialize Inputs
		clk = 0;

		// Wait 100 ns for global reset to finish
		#100;
		clk=1;
        
		// Add stimulus here

	end
   initial forever
	begin
	#1;
	clk=~clk;
	end 
endmodule

